library verilog;
use verilog.vl_types.all;
entity DE2_115 is
    port(
        CLOCK_50        : in     vl_logic;
        CLOCK2_50       : in     vl_logic;
        CLOCK3_50       : in     vl_logic;
        SMA_CLKIN       : in     vl_logic;
        SMA_CLKOUT      : out    vl_logic;
        LEDG            : out    vl_logic_vector(8 downto 0);
        LEDR            : out    vl_logic_vector(17 downto 0);
        KEY             : in     vl_logic_vector(3 downto 0);
        EX_IO           : inout  vl_logic_vector(6 downto 0);
        SW              : in     vl_logic_vector(17 downto 0);
        HEX0            : out    vl_logic_vector(6 downto 0);
        HEX1            : out    vl_logic_vector(6 downto 0);
        HEX2            : out    vl_logic_vector(6 downto 0);
        HEX3            : out    vl_logic_vector(6 downto 0);
        HEX4            : out    vl_logic_vector(6 downto 0);
        HEX5            : out    vl_logic_vector(6 downto 0);
        HEX6            : out    vl_logic_vector(6 downto 0);
        HEX7            : out    vl_logic_vector(6 downto 0);
        LCD_BLON        : out    vl_logic;
        LCD_DATA        : inout  vl_logic_vector(7 downto 0);
        LCD_EN          : out    vl_logic;
        LCD_ON          : out    vl_logic;
        LCD_RS          : out    vl_logic;
        LCD_RW          : out    vl_logic;
        UART_CTS        : in     vl_logic;
        UART_RTS        : out    vl_logic;
        UART_RXD        : in     vl_logic;
        UART_TXD        : out    vl_logic;
        PS2_CLK         : inout  vl_logic;
        PS2_CLK2        : inout  vl_logic;
        PS2_DAT         : inout  vl_logic;
        PS2_DAT2        : inout  vl_logic;
        SD_CLK          : out    vl_logic;
        SD_CMD          : inout  vl_logic;
        SD_DAT          : inout  vl_logic_vector(3 downto 0);
        SD_WP_N         : in     vl_logic;
        VGA_B           : out    vl_logic_vector(7 downto 0);
        VGA_BLANK_N     : out    vl_logic;
        VGA_CLK         : out    vl_logic;
        VGA_G           : out    vl_logic_vector(7 downto 0);
        VGA_HS          : out    vl_logic;
        VGA_R           : out    vl_logic_vector(7 downto 0);
        VGA_SYNC_N      : out    vl_logic;
        VGA_VS          : out    vl_logic;
        AUD_ADCDAT      : in     vl_logic;
        AUD_ADCLRCK     : inout  vl_logic;
        AUD_BCLK        : inout  vl_logic;
        AUD_DACDAT      : out    vl_logic;
        AUD_DACLRCK     : inout  vl_logic;
        AUD_XCK         : out    vl_logic;
        EEP_I2C_SCLK    : out    vl_logic;
        EEP_I2C_SDAT    : inout  vl_logic;
        I2C_SCLK        : out    vl_logic;
        I2C_SDAT        : inout  vl_logic;
        ENET0_GTX_CLK   : out    vl_logic;
        ENET0_INT_N     : in     vl_logic;
        ENET0_LINK100   : in     vl_logic;
        ENET0_MDC       : out    vl_logic;
        ENET0_MDIO      : inout  vl_logic;
        ENET0_RST_N     : out    vl_logic;
        ENET0_RX_CLK    : in     vl_logic;
        ENET0_RX_COL    : in     vl_logic;
        ENET0_RX_CRS    : in     vl_logic;
        ENET0_RX_DATA   : in     vl_logic_vector(3 downto 0);
        ENET0_RX_DV     : in     vl_logic;
        ENET0_RX_ER     : in     vl_logic;
        ENET0_TX_CLK    : in     vl_logic;
        ENET0_TX_DATA   : out    vl_logic_vector(3 downto 0);
        ENET0_TX_EN     : out    vl_logic;
        ENET0_TX_ER     : out    vl_logic;
        ENETCLK_25      : in     vl_logic;
        ENET1_GTX_CLK   : out    vl_logic;
        ENET1_INT_N     : in     vl_logic;
        ENET1_LINK100   : in     vl_logic;
        ENET1_MDC       : out    vl_logic;
        ENET1_MDIO      : inout  vl_logic;
        ENET1_RST_N     : out    vl_logic;
        ENET1_RX_CLK    : in     vl_logic;
        ENET1_RX_COL    : in     vl_logic;
        ENET1_RX_CRS    : in     vl_logic;
        ENET1_RX_DATA   : in     vl_logic_vector(3 downto 0);
        ENET1_RX_DV     : in     vl_logic;
        ENET1_RX_ER     : in     vl_logic;
        ENET1_TX_CLK    : in     vl_logic;
        ENET1_TX_DATA   : out    vl_logic_vector(3 downto 0);
        ENET1_TX_EN     : out    vl_logic;
        ENET1_TX_ER     : out    vl_logic;
        TD_CLK27        : in     vl_logic;
        TD_DATA         : in     vl_logic_vector(7 downto 0);
        TD_HS           : in     vl_logic;
        TD_RESET_N      : out    vl_logic;
        TD_VS           : in     vl_logic;
        OTG_ADDR        : out    vl_logic_vector(1 downto 0);
        OTG_CS_N        : out    vl_logic;
        OTG_DATA        : inout  vl_logic_vector(15 downto 0);
        OTG_INT         : in     vl_logic;
        OTG_RD_N        : out    vl_logic;
        OTG_RST_N       : out    vl_logic;
        OTG_WE_N        : out    vl_logic;
        IRDA_RXD        : in     vl_logic;
        DRAM_ADDR       : out    vl_logic_vector(12 downto 0);
        DRAM_BA         : out    vl_logic_vector(1 downto 0);
        DRAM_CAS_N      : out    vl_logic;
        DRAM_CKE        : out    vl_logic;
        DRAM_CLK        : out    vl_logic;
        DRAM_CS_N       : out    vl_logic;
        DRAM_DQ         : inout  vl_logic_vector(31 downto 0);
        DRAM_DQM        : out    vl_logic_vector(3 downto 0);
        DRAM_RAS_N      : out    vl_logic;
        DRAM_WE_N       : out    vl_logic;
        SRAM_ADDR       : out    vl_logic_vector(19 downto 0);
        SRAM_CE_N       : out    vl_logic;
        SRAM_DQ         : inout  vl_logic_vector(15 downto 0);
        SRAM_LB_N       : out    vl_logic;
        SRAM_OE_N       : out    vl_logic;
        SRAM_UB_N       : out    vl_logic;
        SRAM_WE_N       : out    vl_logic;
        FL_ADDR         : out    vl_logic_vector(22 downto 0);
        FL_CE_N         : out    vl_logic;
        FL_DQ           : inout  vl_logic_vector(7 downto 0);
        FL_OE_N         : out    vl_logic;
        FL_RST_N        : out    vl_logic;
        FL_RY           : in     vl_logic;
        FL_WE_N         : out    vl_logic;
        FL_WP_N         : out    vl_logic
    );
end DE2_115;
