library verilog;
use verilog.vl_types.all;
entity toplevel is
end toplevel;
