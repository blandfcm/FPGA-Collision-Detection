`timescale 1ns / 1ps

module toplevel;

reg CLK = 1'b0;
reg[31:0] p1x;
reg[31:0] p1y;
reg[31:0] p1z;
reg[31:0] p1r;
reg[31:0] p2x;
reg[31:0] p2y;
reg[31:0] p2z;
reg[2:0] s0, s1, s2;
/*wire[31:0] s0, s1;
	assign s0 = 32'b01000000100000000000000000000000;
	assign s1 = 32'b01000000000000000000000000000000;
*/
//reg[31:0] s2;
reg[31:0] R9, R10;
reg[31:0] g1c, g2c;
wire[31:0] cX, cY, cZ, nx, ny, nz, depthC;
	assign cX = 32'b10111111001101110110010000000110; 	//-0.71637
	assign cY = 32'b10111110110101100100011110011001; 	//-0.418515
	assign cZ = 32'b00111111000011101110101001100100; 	//0.558264
	assign nx = 32'b10111110011000110011011100100010; 	//-0.22189
	assign ny = 32'b10111111000111110011011011011111; 	//-0.621931
	assign nz = 32'b10111111010000000100000000000111; 	//-0.750977
	assign depthC = 32'b00111111001010010101011111011110; 	//0.661497
wire[31:0] check;
wire ret_val, done_flag;
reg rst_wire;

dCollideSphereBox test0(
	.rst(rst_wire),
	.clk(CLK),
	.x1(p1x), 	
	.y1(p1y), 	
	.z1(p1z), 	
	.x2(p2x), 	
	.y2(p2y), 	
	.z2(p2z),	
	//.side0(s0),
	//.side1(s1),
	//.side2(s2),
	.r0(cX),
	.r1(cY),
	.r2(cZ),
	.r4(nx),
	.r5(ny),
	.r6(nz),
	.r8(depthC),
	//.r9(s0),
	//.r10(s1),
	//.side2(s2),
	.r9(R9),
	.r10(R10),
	/*.cx(cX), 
	.cy(cY), 
	.cz(cZ),
	.normalx(nx), 
	.normaly(ny), 
	.normalz(nz),
	.depth(depthC),*/
	.ret(ret_val), 
	.done(done_flag)
);


integer i;

initial
begin
CLK = 0;
rst_wire = 0;
	p1x = 32'b11000001100011111011000010011010; 	//-17.961231
	p1y = 32'b10111111000101001100011100011001; 	//-0.581163
	p1z = 32'b01000000111111100101101101101110; 	//7.948661
	p2x = 32'b11000001100000011101100011010010; 	//-16.23087
	p2y = 32'b00111111101001110100011010110010; 	//1.306845
	p2z = 32'b01000001000101001110100110110011;	//9.307055
	//s0 = 3'd4;
	//s1 = 3'd2;
	//s2 = 3'd0;
	/*s0 = 32'b01000000100000000000000000000000;	//4.0
	s1 = 32'b01000000000000000000000000000000;	//2.0
	s2 = 32'b00111111100000000000000000000000;	//1.0*/
	
	R9 = 32'b10111111001010010110111100010001; 	//-0.661851
	R10 = 32'b00111110101101001001000100001000; 	//0.352669
end

always  
    #1  CLK =  ! CLK; 
initial 
	#10000  $stop; 

endmodule