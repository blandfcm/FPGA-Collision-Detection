library verilog;
use verilog.vl_types.all;
entity toplevel0 is
end toplevel0;
