module dCollideSpheres(x1, y1, z1, r1, x2, y2, z2, r2, cx, cy, cz, normalX, normalY, normalZ, depth, g1, g2, return);
/**
	dVector3 p1:		x1, y1, z1
	dReal r1:			r1
	dVector3 p2:		x2, y2, z2
	dReal r2:			r2
	dContactGeom *c:	
		dVector3 pos		cx, cy, cz
		dVector3 normal	normalX, normalY, normalZ
		dReal depth			depth
		dGeomID g1, g2		g1, g2
*/
