module Collision_Detection();

endmodule
